module porta_or
(
	input a, b,
	output s
);

	assign s = a | b;

endmodule 