module porta_and
(
	input a, b,
	output s
);

	assign s = a & b;
	
endmodule 