module igualdade_complemento_1
(
	input A, M,
	output S
);

	assign S = A ^ M;
	
endmodule 